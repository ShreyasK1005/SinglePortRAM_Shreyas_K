package ram_package;
// `include "ram_package.sv"
 `include "ram_transaction.sv"
 `include "ram_generator.sv"
 `include "ram_driver.sv"
 `include "ram_monitor.sv"
 `include "ram_reference_model.sv"
 `include "ram_scoreboard.sv"
 `include "ram_environment.sv"
 `include "ram_test.sv"
endpackage